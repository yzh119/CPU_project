`include "macros.v"

module hi_lo_reg (
	
);

endmodule